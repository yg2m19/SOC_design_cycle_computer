// Example code for an M0 AHBLite System
//  Iain McNally
//  ECS, University of Soutampton
//
// This module is an AHB-Lite Slave containing a ROM
//
// Number of addressable locations : 2**MEMWIDTH
// Size of each addressable location : 8 bits
// Supported transfer sizes : Word, Halfword, Byte
// Alignment of base address : Word aligned
//

`define STRINGIFY(x) `"x`"

`ifdef prog_file
  // already defined - do nothing
`else
  `define prog_file  code.hex
`endif

module ahb_rom #(
  parameter MEMWIDTH = 14
)(
  //AHBLITE INTERFACE

    //Slave Select Signal
    input HSEL,
    //Global Signals
    input HCLK,
    input HRESETn,
    //Address, Control & Write Data
    input HREADY,
    input [31:0] HADDR,
    input [1:0] HTRANS,
    input HWRITE,
    input [2:0] HSIZE,
    input [31:0] HWDATA,
    // Transfer Response & Read Data
    output HREADYOUT,
    output [31:0] HRDATA

);

timeunit 1ns;
timeprecision 100ps;

  localparam No_Transfer = 2'b0;

// Memory Array  
  logic [31:0] memory[0:(2**(MEMWIDTH-2)-1)];

//control signals are stored in registers
  logic read_enable;
  logic [MEMWIDTH-2:0] word_address;
  logic [3:0] byte_select;
  

// read program from "code.hex" rom

  assign memory[ 0 ] = 32'h20000100;
  assign memory[ 1 ] = 32'h000000C1;
  assign memory[ 2 ] = 32'h000000ED;
  assign memory[ 3 ] = 32'h000000F1;
  assign memory[ 4 ] = 32'h000000F5;
  assign memory[ 5 ] = 32'h000000F9;
  assign memory[ 6 ] = 32'h000000FD;
  assign memory[ 7 ] = 32'h00000000;
  assign memory[ 8 ] = 32'h00000000;
  assign memory[ 9 ] = 32'h00000000;
  assign memory[ 10 ] = 32'h00000000;
  assign memory[ 11 ] = 32'h00000101;
  assign memory[ 12 ] = 32'h00000105;
  assign memory[ 13 ] = 32'h00000000;
  assign memory[ 14 ] = 32'h00000109;
  assign memory[ 15 ] = 32'h0000010D;
  assign memory[ 16 ] = 32'h00000111;
  assign memory[ 17 ] = 32'h00000111;
  assign memory[ 18 ] = 32'h00000111;
  assign memory[ 19 ] = 32'h00000111;
  assign memory[ 20 ] = 32'h00000111;
  assign memory[ 21 ] = 32'h00000111;
  assign memory[ 22 ] = 32'h00000111;
  assign memory[ 23 ] = 32'h00000111;
  assign memory[ 24 ] = 32'h00000111;
  assign memory[ 25 ] = 32'h00000111;
  assign memory[ 26 ] = 32'h00000111;
  assign memory[ 27 ] = 32'h00000111;
  assign memory[ 28 ] = 32'h00000111;
  assign memory[ 29 ] = 32'h00000115;
  assign memory[ 30 ] = 32'h00000119;
  assign memory[ 31 ] = 32'h0000011D;
  assign memory[ 32 ] = 32'h00000121;
  assign memory[ 33 ] = 32'h00000125;
  assign memory[ 34 ] = 32'h00000129;
  assign memory[ 35 ] = 32'h0000012D;
  assign memory[ 36 ] = 32'h00000131;
  assign memory[ 37 ] = 32'h00000135;
  assign memory[ 38 ] = 32'h00000000;
  assign memory[ 39 ] = 32'h00000000;
  assign memory[ 40 ] = 32'h00000139;
  assign memory[ 41 ] = 32'h0000013D;
  assign memory[ 42 ] = 32'h00000141;
  assign memory[ 43 ] = 32'h00000000;
  assign memory[ 44 ] = 32'h00000145;
  assign memory[ 45 ] = 32'h00000149;
  assign memory[ 46 ] = 32'h0000014D;
  assign memory[ 47 ] = 32'h00000151;
  assign memory[ 48 ] = 32'hB083B500;
  assign memory[ 49 ] = 32'h93014B07;
  assign memory[ 50 ] = 32'h9B01E004;
  assign memory[ 51 ] = 32'h92011D1A;
  assign memory[ 52 ] = 32'h601A2200;
  assign memory[ 53 ] = 32'h4B049A01;
  assign memory[ 54 ] = 32'hD3F6429A;
  assign memory[ 55 ] = 32'hF922F000;
  assign memory[ 56 ] = 32'h46C0E7FE;
  assign memory[ 57 ] = 32'h20000000;
  assign memory[ 58 ] = 32'h20000000;
  assign memory[ 59 ] = 32'h46C0E7FE;
  assign memory[ 60 ] = 32'h46C0E7FE;
  assign memory[ 61 ] = 32'h46C0E7FE;
  assign memory[ 62 ] = 32'h46C0E7FE;
  assign memory[ 63 ] = 32'h46C0E7FE;
  assign memory[ 64 ] = 32'h46C0E7FE;
  assign memory[ 65 ] = 32'h46C0E7FE;
  assign memory[ 66 ] = 32'h46C0E7FE;
  assign memory[ 67 ] = 32'h46C0E7FE;
  assign memory[ 68 ] = 32'h46C0E7FE;
  assign memory[ 69 ] = 32'h46C0E7FE;
  assign memory[ 70 ] = 32'h46C0E7FE;
  assign memory[ 71 ] = 32'h46C0E7FE;
  assign memory[ 72 ] = 32'h46C0E7FE;
  assign memory[ 73 ] = 32'h46C0E7FE;
  assign memory[ 74 ] = 32'h46C0E7FE;
  assign memory[ 75 ] = 32'h46C0E7FE;
  assign memory[ 76 ] = 32'h46C0E7FE;
  assign memory[ 77 ] = 32'h46C0E7FE;
  assign memory[ 78 ] = 32'h46C0E7FE;
  assign memory[ 79 ] = 32'h46C0E7FE;
  assign memory[ 80 ] = 32'h46C0E7FE;
  assign memory[ 81 ] = 32'h46C0E7FE;
  assign memory[ 82 ] = 32'h46C0E7FE;
  assign memory[ 83 ] = 32'h46C0E7FE;
  assign memory[ 84 ] = 32'h46C0E7FE;
  assign memory[ 85 ] = 32'h9001B082;
  assign memory[ 86 ] = 32'h681B4B05;
  assign memory[ 87 ] = 32'h22013304;
  assign memory[ 88 ] = 32'h4B03601A;
  assign memory[ 89 ] = 32'h9A01681B;
  assign memory[ 90 ] = 32'h46C0601A;
  assign memory[ 91 ] = 32'h4770B002;
  assign memory[ 92 ] = 32'h0000117C;
  assign memory[ 93 ] = 32'h681B4B02;
  assign memory[ 94 ] = 32'h0018681B;
  assign memory[ 95 ] = 32'h46C04770;
  assign memory[ 96 ] = 32'h0000117C;
  assign memory[ 97 ] = 32'h9001B082;
  assign memory[ 98 ] = 32'h681A4B04;
  assign memory[ 99 ] = 32'h009B9B01;
  assign memory[ 100 ] = 32'h681B18D3;
  assign memory[ 101 ] = 32'hB0020018;
  assign memory[ 102 ] = 32'h46C04770;
  assign memory[ 103 ] = 32'h00001178;
  assign memory[ 104 ] = 32'h2314B082;
  assign memory[ 105 ] = 32'hE00B9301;
  assign memory[ 106 ] = 32'h93002323;
  assign memory[ 107 ] = 32'h9B00E002;
  assign memory[ 108 ] = 32'h93003B01;
  assign memory[ 109 ] = 32'h2B009B00;
  assign memory[ 110 ] = 32'h9B01DCF9;
  assign memory[ 111 ] = 32'h93013B01;
  assign memory[ 112 ] = 32'h2B009B01;
  assign memory[ 113 ] = 32'h46C0DCF0;
  assign memory[ 114 ] = 32'h4770B002;
  assign memory[ 115 ] = 32'hB085B500;
  assign memory[ 116 ] = 32'h91009001;
  assign memory[ 117 ] = 32'h9A009B01;
  assign memory[ 118 ] = 32'h0013435A;
  assign memory[ 119 ] = 32'h189B009B;
  assign memory[ 120 ] = 32'h4908005B;
  assign memory[ 121 ] = 32'hF0000018;
  assign memory[ 122 ] = 32'h0003FE7F;
  assign memory[ 123 ] = 32'h9B039303;
  assign memory[ 124 ] = 32'h05D22280;
  assign memory[ 125 ] = 32'h44634694;
  assign memory[ 126 ] = 32'h9B029302;
  assign memory[ 127 ] = 32'hB0050018;
  assign memory[ 128 ] = 32'h46C0BD00;
  assign memory[ 129 ] = 32'h000F4240;
  assign memory[ 130 ] = 32'hB087B500;
  assign memory[ 131 ] = 32'h9B019001;
  assign memory[ 132 ] = 32'h00184910;
  assign memory[ 133 ] = 32'hFE68F000;
  assign memory[ 134 ] = 32'h93050003;
  assign memory[ 135 ] = 32'h4A0E9B05;
  assign memory[ 136 ] = 32'h9B01435A;
  assign memory[ 137 ] = 32'h490D18D3;
  assign memory[ 138 ] = 32'hF0000018;
  assign memory[ 139 ] = 32'h0003FE5D;
  assign memory[ 140 ] = 32'h9B059304;
  assign memory[ 141 ] = 32'h435A2264;
  assign memory[ 142 ] = 32'h18D39B04;
  assign memory[ 143 ] = 32'h9B039303;
  assign memory[ 144 ] = 32'h05D222C0;
  assign memory[ 145 ] = 32'h44634694;
  assign memory[ 146 ] = 32'h9B029302;
  assign memory[ 147 ] = 32'hB0070018;
  assign memory[ 148 ] = 32'h46C0BD00;
  assign memory[ 149 ] = 32'h02BF2000;
  assign memory[ 150 ] = 32'hFD40E000;
  assign memory[ 151 ] = 32'h000BB800;
  assign memory[ 152 ] = 32'hB085B500;
  assign memory[ 153 ] = 32'h99019001;
  assign memory[ 154 ] = 32'hF000480B;
  assign memory[ 155 ] = 32'h1E03FE3D;
  assign memory[ 156 ] = 32'h2380D102;
  assign memory[ 157 ] = 32'hE00C061B;
  assign memory[ 158 ] = 32'h48079901;
  assign memory[ 159 ] = 32'hFE34F000;
  assign memory[ 160 ] = 32'h93030003;
  assign memory[ 161 ] = 32'h22809B03;
  assign memory[ 162 ] = 32'h46940612;
  assign memory[ 163 ] = 32'h93024463;
  assign memory[ 164 ] = 32'h00189B02;
  assign memory[ 165 ] = 32'hBD00B005;
  assign memory[ 166 ] = 32'h000BB800;
  assign memory[ 167 ] = 32'hB089B500;
  assign memory[ 168 ] = 32'h91009001;
  assign memory[ 169 ] = 32'h2B009B01;
  assign memory[ 170 ] = 32'h2300D104;
  assign memory[ 171 ] = 32'h23009307;
  assign memory[ 172 ] = 32'hE01B9306;
  assign memory[ 173 ] = 32'h48179901;
  assign memory[ 174 ] = 32'hFE16F000;
  assign memory[ 175 ] = 32'h93050003;
  assign memory[ 176 ] = 32'h9A059B00;
  assign memory[ 177 ] = 32'h49144353;
  assign memory[ 178 ] = 32'hF0000018;
  assign memory[ 179 ] = 32'h0003FE0D;
  assign memory[ 180 ] = 32'h9B009307;
  assign memory[ 181 ] = 32'h435A9A05;
  assign memory[ 182 ] = 32'h49109B07;
  assign memory[ 183 ] = 32'h18D3434B;
  assign memory[ 184 ] = 32'h0018490F;
  assign memory[ 185 ] = 32'hFE00F000;
  assign memory[ 186 ] = 32'h93060003;
  assign memory[ 187 ] = 32'h00139A07;
  assign memory[ 188 ] = 32'h189B009B;
  assign memory[ 189 ] = 32'h001A005B;
  assign memory[ 190 ] = 32'h18D39B06;
  assign memory[ 191 ] = 32'h9B049304;
  assign memory[ 192 ] = 32'h061222A0;
  assign memory[ 193 ] = 32'h44634694;
  assign memory[ 194 ] = 32'h9B039303;
  assign memory[ 195 ] = 32'hB0090018;
  assign memory[ 196 ] = 32'h46C0BD00;
  assign memory[ 197 ] = 32'h1B774000;
  assign memory[ 198 ] = 32'h00989680;
  assign memory[ 199 ] = 32'hFF676980;
  assign memory[ 200 ] = 32'h000F4240;
  assign memory[ 201 ] = 32'hB096B510;
  assign memory[ 202 ] = 32'h93152300;
  assign memory[ 203 ] = 32'h93142300;
  assign memory[ 204 ] = 32'h93102300;
  assign memory[ 205 ] = 32'h93112300;
  assign memory[ 206 ] = 32'h930E2300;
  assign memory[ 207 ] = 32'h930F2300;
  assign memory[ 208 ] = 32'h930D2300;
  assign memory[ 209 ] = 32'h93082300;
  assign memory[ 210 ] = 32'h93072300;
  assign memory[ 211 ] = 32'h93062300;
  assign memory[ 212 ] = 32'h93052300;
  assign memory[ 213 ] = 32'h93042300;
  assign memory[ 214 ] = 32'h93032300;
  assign memory[ 215 ] = 32'h93134BDA;
  assign memory[ 216 ] = 32'h93122300;
  assign memory[ 217 ] = 32'h93022300;
  assign memory[ 218 ] = 32'h930C2306;
  assign memory[ 219 ] = 32'h930B2303;
  assign memory[ 220 ] = 32'h930A2301;
  assign memory[ 221 ] = 32'h93092302;
  assign memory[ 222 ] = 32'h93012300;
  assign memory[ 223 ] = 32'hF7FF2000;
  assign memory[ 224 ] = 32'h0003FF01;
  assign memory[ 225 ] = 32'h20019308;
  assign memory[ 226 ] = 32'hFEFCF7FF;
  assign memory[ 227 ] = 32'h93070003;
  assign memory[ 228 ] = 32'hF7FF2005;
  assign memory[ 229 ] = 32'h0003FEF7;
  assign memory[ 230 ] = 32'h9A139303;
  assign memory[ 231 ] = 32'h00119B03;
  assign memory[ 232 ] = 32'hF7FF0018;
  assign memory[ 233 ] = 32'h0003FF7B;
  assign memory[ 234 ] = 32'h9B029302;
  assign memory[ 235 ] = 32'h05D222C0;
  assign memory[ 236 ] = 32'h44634694;
  assign memory[ 237 ] = 32'h9A019301;
  assign memory[ 238 ] = 32'h429A9B12;
  assign memory[ 239 ] = 32'h9B01DD01;
  assign memory[ 240 ] = 32'h9A079312;
  assign memory[ 241 ] = 32'h005B23A0;
  assign memory[ 242 ] = 32'hDD06429A;
  assign memory[ 243 ] = 32'h23A09A08;
  assign memory[ 244 ] = 32'h429A005B;
  assign memory[ 245 ] = 32'h2301DD01;
  assign memory[ 246 ] = 32'h9B07930D;
  assign memory[ 247 ] = 32'hD1182B00;
  assign memory[ 248 ] = 32'h2B009B08;
  assign memory[ 249 ] = 32'h9B0DD115;
  assign memory[ 250 ] = 32'hD1122B01;
  assign memory[ 251 ] = 32'h93142301;
  assign memory[ 252 ] = 32'h93112303;
  assign memory[ 253 ] = 32'h930D2300;
  assign memory[ 254 ] = 32'h930F2300;
  assign memory[ 255 ] = 32'h930E2300;
  assign memory[ 256 ] = 32'hF7FF2000;
  assign memory[ 257 ] = 32'hF7FFFEA7;
  assign memory[ 258 ] = 32'h4BB0FECB;
  assign memory[ 259 ] = 32'hF7FF0018;
  assign memory[ 260 ] = 32'h9B14FEA1;
  assign memory[ 261 ] = 32'hD1012B00;
  assign memory[ 262 ] = 32'hFCC3F000;
  assign memory[ 263 ] = 32'h23409A08;
  assign memory[ 264 ] = 32'h429A33FF;
  assign memory[ 265 ] = 32'h9B07DD04;
  assign memory[ 266 ] = 32'hD1012B00;
  assign memory[ 267 ] = 32'h930E2301;
  assign memory[ 268 ] = 32'h2B009B08;
  assign memory[ 269 ] = 32'h9B0ED110;
  assign memory[ 270 ] = 32'hD10D2B01;
  assign memory[ 271 ] = 32'h2B009B07;
  assign memory[ 272 ] = 32'h9B10D10A;
  assign memory[ 273 ] = 32'hDC032B08;
  assign memory[ 274 ] = 32'h33019B10;
  assign memory[ 275 ] = 32'hE0019310;
  assign memory[ 276 ] = 32'h93102300;
  assign memory[ 277 ] = 32'h930E2300;
  assign memory[ 278 ] = 32'h23409A07;
  assign memory[ 279 ] = 32'h429A33FF;
  assign memory[ 280 ] = 32'h9B08DD04;
  assign memory[ 281 ] = 32'hD1012B00;
  assign memory[ 282 ] = 32'h930F2301;
  assign memory[ 283 ] = 32'h2B009B07;
  assign memory[ 284 ] = 32'h9B0FD13E;
  assign memory[ 285 ] = 32'hD13B2B01;
  assign memory[ 286 ] = 32'h2B009B08;
  assign memory[ 287 ] = 32'h9B11D138;
  assign memory[ 288 ] = 32'hDD072B00;
  assign memory[ 289 ] = 32'h3B019B11;
  assign memory[ 290 ] = 32'h23009311;
  assign memory[ 291 ] = 32'h23009310;
  assign memory[ 292 ] = 32'hE02D930F;
  assign memory[ 293 ] = 32'h22FA9B09;
  assign memory[ 294 ] = 32'h435A0092;
  assign memory[ 295 ] = 32'h21649B0A;
  assign memory[ 296 ] = 32'h18D1434B;
  assign memory[ 297 ] = 32'h00139A0B;
  assign memory[ 298 ] = 32'h189B009B;
  assign memory[ 299 ] = 32'h18CA005B;
  assign memory[ 300 ] = 32'h18D39B0C;
  assign memory[ 301 ] = 32'h23009313;
  assign memory[ 302 ] = 32'h23009314;
  assign memory[ 303 ] = 32'h23009315;
  assign memory[ 304 ] = 32'h9B09930F;
  assign memory[ 305 ] = 32'h009222FA;
  assign memory[ 306 ] = 32'h9B0A435A;
  assign memory[ 307 ] = 32'h434B2164;
  assign memory[ 308 ] = 32'h9A0B18D1;
  assign memory[ 309 ] = 32'h009B0013;
  assign memory[ 310 ] = 32'h005B189B;
  assign memory[ 311 ] = 32'h9B0C18CA;
  assign memory[ 312 ] = 32'h228018D3;
  assign memory[ 313 ] = 32'h46940592;
  assign memory[ 314 ] = 32'h00184463;
  assign memory[ 315 ] = 32'hFE32F7FF;
  assign memory[ 316 ] = 32'h2B019B11;
  assign memory[ 317 ] = 32'hE122D100;
  assign memory[ 318 ] = 32'h2B00DC03;
  assign memory[ 319 ] = 32'hF000D009;
  assign memory[ 320 ] = 32'h2B02FCE9;
  assign memory[ 321 ] = 32'hE229D100;
  assign memory[ 322 ] = 32'hD1002B03;
  assign memory[ 323 ] = 32'hF000E339;
  assign memory[ 324 ] = 32'h9B10FCE1;
  assign memory[ 325 ] = 32'hD9012B09;
  assign memory[ 326 ] = 32'hFCD2F000;
  assign memory[ 327 ] = 32'h009A9B10;
  assign memory[ 328 ] = 32'h18D34B6B;
  assign memory[ 329 ] = 32'h469F681B;
  assign memory[ 330 ] = 32'h930C2300;
  assign memory[ 331 ] = 32'h22FA9B09;
  assign memory[ 332 ] = 32'h435A0092;
  assign memory[ 333 ] = 32'h21649B0A;
  assign memory[ 334 ] = 32'h18D1434B;
  assign memory[ 335 ] = 32'h00139A0B;
  assign memory[ 336 ] = 32'h189B009B;
  assign memory[ 337 ] = 32'h18CA005B;
  assign memory[ 338 ] = 32'h18D39B0C;
  assign memory[ 339 ] = 32'h05922280;
  assign memory[ 340 ] = 32'h44634694;
  assign memory[ 341 ] = 32'hF7FF0018;
  assign memory[ 342 ] = 32'hE0EFFDFD;
  assign memory[ 343 ] = 32'h930C2301;
  assign memory[ 344 ] = 32'h22FA9B09;
  assign memory[ 345 ] = 32'h435A0092;
  assign memory[ 346 ] = 32'h21649B0A;
  assign memory[ 347 ] = 32'h18D1434B;
  assign memory[ 348 ] = 32'h00139A0B;
  assign memory[ 349 ] = 32'h189B009B;
  assign memory[ 350 ] = 32'h18CA005B;
  assign memory[ 351 ] = 32'h18D39B0C;
  assign memory[ 352 ] = 32'h05922280;
  assign memory[ 353 ] = 32'h44634694;
  assign memory[ 354 ] = 32'hF7FF0018;
  assign memory[ 355 ] = 32'hE0D5FDE3;
  assign memory[ 356 ] = 32'h930C2302;
  assign memory[ 357 ] = 32'h22FA9B09;
  assign memory[ 358 ] = 32'h435A0092;
  assign memory[ 359 ] = 32'h21649B0A;
  assign memory[ 360 ] = 32'h18D1434B;
  assign memory[ 361 ] = 32'h00139A0B;
  assign memory[ 362 ] = 32'h189B009B;
  assign memory[ 363 ] = 32'h18CA005B;
  assign memory[ 364 ] = 32'h18D39B0C;
  assign memory[ 365 ] = 32'h05922280;
  assign memory[ 366 ] = 32'h44634694;
  assign memory[ 367 ] = 32'hF7FF0018;
  assign memory[ 368 ] = 32'hE0BBFDC9;
  assign memory[ 369 ] = 32'h930C2303;
  assign memory[ 370 ] = 32'h22FA9B09;
  assign memory[ 371 ] = 32'h435A0092;
  assign memory[ 372 ] = 32'h21649B0A;
  assign memory[ 373 ] = 32'h18D1434B;
  assign memory[ 374 ] = 32'h00139A0B;
  assign memory[ 375 ] = 32'h189B009B;
  assign memory[ 376 ] = 32'h18CA005B;
  assign memory[ 377 ] = 32'h18D39B0C;
  assign memory[ 378 ] = 32'h05922280;
  assign memory[ 379 ] = 32'h44634694;
  assign memory[ 380 ] = 32'hF7FF0018;
  assign memory[ 381 ] = 32'hE0A1FDAF;
  assign memory[ 382 ] = 32'h930C2304;
  assign memory[ 383 ] = 32'h22FA9B09;
  assign memory[ 384 ] = 32'h435A0092;
  assign memory[ 385 ] = 32'h21649B0A;
  assign memory[ 386 ] = 32'h18D1434B;
  assign memory[ 387 ] = 32'h00139A0B;
  assign memory[ 388 ] = 32'h189B009B;
  assign memory[ 389 ] = 32'h18CA005B;
  assign memory[ 390 ] = 32'h18D39B0C;
  assign memory[ 391 ] = 32'h05922280;
  assign memory[ 392 ] = 32'h44634694;
  assign memory[ 393 ] = 32'hF7FF0018;
  assign memory[ 394 ] = 32'hE087FD95;
  assign memory[ 395 ] = 32'h930C2305;
  assign memory[ 396 ] = 32'h22FA9B09;
  assign memory[ 397 ] = 32'h435A0092;
  assign memory[ 398 ] = 32'h21649B0A;
  assign memory[ 399 ] = 32'h18D1434B;
  assign memory[ 400 ] = 32'h00139A0B;
  assign memory[ 401 ] = 32'h189B009B;
  assign memory[ 402 ] = 32'h18CA005B;
  assign memory[ 403 ] = 32'h18D39B0C;
  assign memory[ 404 ] = 32'h05922280;
  assign memory[ 405 ] = 32'h44634694;
  assign memory[ 406 ] = 32'hF7FF0018;
  assign memory[ 407 ] = 32'hE06DFD7B;
  assign memory[ 408 ] = 32'h930C2306;
  assign memory[ 409 ] = 32'h22FA9B09;
  assign memory[ 410 ] = 32'h435A0092;
  assign memory[ 411 ] = 32'h21649B0A;
  assign memory[ 412 ] = 32'h18D1434B;
  assign memory[ 413 ] = 32'h00139A0B;
  assign memory[ 414 ] = 32'h189B009B;
  assign memory[ 415 ] = 32'h18CA005B;
  assign memory[ 416 ] = 32'h18D39B0C;
  assign memory[ 417 ] = 32'h05922280;
  assign memory[ 418 ] = 32'h44634694;
  assign memory[ 419 ] = 32'hF7FF0018;
  assign memory[ 420 ] = 32'hE053FD61;
  assign memory[ 421 ] = 32'h930C2307;
  assign memory[ 422 ] = 32'h22FA9B09;
  assign memory[ 423 ] = 32'h435A0092;
  assign memory[ 424 ] = 32'h21649B0A;
  assign memory[ 425 ] = 32'h18D1434B;
  assign memory[ 426 ] = 32'h00139A0B;
  assign memory[ 427 ] = 32'h189B009B;
  assign memory[ 428 ] = 32'h18CA005B;
  assign memory[ 429 ] = 32'h18D39B0C;
  assign memory[ 430 ] = 32'h05922280;
  assign memory[ 431 ] = 32'h44634694;
  assign memory[ 432 ] = 32'hF7FF0018;
  assign memory[ 433 ] = 32'hE039FD47;
  assign memory[ 434 ] = 32'h00000858;
  assign memory[ 435 ] = 32'h20000858;
  assign memory[ 436 ] = 32'h000010C0;
  assign memory[ 437 ] = 32'h930C2308;
  assign memory[ 438 ] = 32'h22FA9B09;
  assign memory[ 439 ] = 32'h435A0092;
  assign memory[ 440 ] = 32'h21649B0A;
  assign memory[ 441 ] = 32'h18D1434B;
  assign memory[ 442 ] = 32'h00139A0B;
  assign memory[ 443 ] = 32'h189B009B;
  assign memory[ 444 ] = 32'h18CA005B;
  assign memory[ 445 ] = 32'h18D39B0C;
  assign memory[ 446 ] = 32'h05922280;
  assign memory[ 447 ] = 32'h44634694;
  assign memory[ 448 ] = 32'hF7FF0018;
  assign memory[ 449 ] = 32'hE019FD27;
  assign memory[ 450 ] = 32'h930C2309;
  assign memory[ 451 ] = 32'h22FA9B09;
  assign memory[ 452 ] = 32'h435A0092;
  assign memory[ 453 ] = 32'h21649B0A;
  assign memory[ 454 ] = 32'h18D1434B;
  assign memory[ 455 ] = 32'h00139A0B;
  assign memory[ 456 ] = 32'h189B009B;
  assign memory[ 457 ] = 32'h18CA005B;
  assign memory[ 458 ] = 32'h18D39B0C;
  assign memory[ 459 ] = 32'h05922280;
  assign memory[ 460 ] = 32'h44634694;
  assign memory[ 461 ] = 32'hF7FF0018;
  assign memory[ 462 ] = 32'h46C0FD0D;
  assign memory[ 463 ] = 32'h9B10E3C0;
  assign memory[ 464 ] = 32'hD9002B09;
  assign memory[ 465 ] = 32'h9B10E3BF;
  assign memory[ 466 ] = 32'h4BF1009A;
  assign memory[ 467 ] = 32'h681B18D3;
  assign memory[ 468 ] = 32'h2300469F;
  assign memory[ 469 ] = 32'h9B09930B;
  assign memory[ 470 ] = 32'h009222FA;
  assign memory[ 471 ] = 32'h9B0A435A;
  assign memory[ 472 ] = 32'h434B2164;
  assign memory[ 473 ] = 32'h9A0B18D1;
  assign memory[ 474 ] = 32'h009B0013;
  assign memory[ 475 ] = 32'h005B189B;
  assign memory[ 476 ] = 32'h9B0C18CA;
  assign memory[ 477 ] = 32'h228018D3;
  assign memory[ 478 ] = 32'h46940592;
  assign memory[ 479 ] = 32'h00184463;
  assign memory[ 480 ] = 32'hFCE8F7FF;
  assign memory[ 481 ] = 32'h2301E0E9;
  assign memory[ 482 ] = 32'h9B09930B;
  assign memory[ 483 ] = 32'h009222FA;
  assign memory[ 484 ] = 32'h9B0A435A;
  assign memory[ 485 ] = 32'h434B2164;
  assign memory[ 486 ] = 32'h9A0B18D1;
  assign memory[ 487 ] = 32'h009B0013;
  assign memory[ 488 ] = 32'h005B189B;
  assign memory[ 489 ] = 32'h9B0C18CA;
  assign memory[ 490 ] = 32'h228018D3;
  assign memory[ 491 ] = 32'h46940592;
  assign memory[ 492 ] = 32'h00184463;
  assign memory[ 493 ] = 32'hFCCEF7FF;
  assign memory[ 494 ] = 32'h2302E0CF;
  assign memory[ 495 ] = 32'h9B09930B;
  assign memory[ 496 ] = 32'h009222FA;
  assign memory[ 497 ] = 32'h9B0A435A;
  assign memory[ 498 ] = 32'h434B2164;
  assign memory[ 499 ] = 32'h9A0B18D1;
  assign memory[ 500 ] = 32'h009B0013;
  assign memory[ 501 ] = 32'h005B189B;
  assign memory[ 502 ] = 32'h9B0C18CA;
  assign memory[ 503 ] = 32'h228018D3;
  assign memory[ 504 ] = 32'h46940592;
  assign memory[ 505 ] = 32'h00184463;
  assign memory[ 506 ] = 32'hFCB4F7FF;
  assign memory[ 507 ] = 32'h2303E0B5;
  assign memory[ 508 ] = 32'h9B09930B;
  assign memory[ 509 ] = 32'h009222FA;
  assign memory[ 510 ] = 32'h9B0A435A;
  assign memory[ 511 ] = 32'h434B2164;
  assign memory[ 512 ] = 32'h9A0B18D1;
  assign memory[ 513 ] = 32'h009B0013;
  assign memory[ 514 ] = 32'h005B189B;
  assign memory[ 515 ] = 32'h9B0C18CA;
  assign memory[ 516 ] = 32'h228018D3;
  assign memory[ 517 ] = 32'h46940592;
  assign memory[ 518 ] = 32'h00184463;
  assign memory[ 519 ] = 32'hFC9AF7FF;
  assign memory[ 520 ] = 32'h2304E09B;
  assign memory[ 521 ] = 32'h9B09930B;
  assign memory[ 522 ] = 32'h009222FA;
  assign memory[ 523 ] = 32'h9B0A435A;
  assign memory[ 524 ] = 32'h434B2164;
  assign memory[ 525 ] = 32'h9A0B18D1;
  assign memory[ 526 ] = 32'h009B0013;
  assign memory[ 527 ] = 32'h005B189B;
  assign memory[ 528 ] = 32'h9B0C18CA;
  assign memory[ 529 ] = 32'h228018D3;
  assign memory[ 530 ] = 32'h46940592;
  assign memory[ 531 ] = 32'h00184463;
  assign memory[ 532 ] = 32'hFC80F7FF;
  assign memory[ 533 ] = 32'h2305E081;
  assign memory[ 534 ] = 32'h9B09930B;
  assign memory[ 535 ] = 32'h009222FA;
  assign memory[ 536 ] = 32'h9B0A435A;
  assign memory[ 537 ] = 32'h434B2164;
  assign memory[ 538 ] = 32'h9A0B18D1;
  assign memory[ 539 ] = 32'h009B0013;
  assign memory[ 540 ] = 32'h005B189B;
  assign memory[ 541 ] = 32'h9B0C18CA;
  assign memory[ 542 ] = 32'h228018D3;
  assign memory[ 543 ] = 32'h46940592;
  assign memory[ 544 ] = 32'h00184463;
  assign memory[ 545 ] = 32'hFC66F7FF;
  assign memory[ 546 ] = 32'h2306E067;
  assign memory[ 547 ] = 32'h9B09930B;
  assign memory[ 548 ] = 32'h009222FA;
  assign memory[ 549 ] = 32'h9B0A435A;
  assign memory[ 550 ] = 32'h434B2164;
  assign memory[ 551 ] = 32'h9A0B18D1;
  assign memory[ 552 ] = 32'h009B0013;
  assign memory[ 553 ] = 32'h005B189B;
  assign memory[ 554 ] = 32'h9B0C18CA;
  assign memory[ 555 ] = 32'h228018D3;
  assign memory[ 556 ] = 32'h46940592;
  assign memory[ 557 ] = 32'h00184463;
  assign memory[ 558 ] = 32'hFC4CF7FF;
  assign memory[ 559 ] = 32'h2307E04D;
  assign memory[ 560 ] = 32'h9B09930B;
  assign memory[ 561 ] = 32'h009222FA;
  assign memory[ 562 ] = 32'h9B0A435A;
  assign memory[ 563 ] = 32'h434B2164;
  assign memory[ 564 ] = 32'h9A0B18D1;
  assign memory[ 565 ] = 32'h009B0013;
  assign memory[ 566 ] = 32'h005B189B;
  assign memory[ 567 ] = 32'h9B0C18CA;
  assign memory[ 568 ] = 32'h228018D3;
  assign memory[ 569 ] = 32'h46940592;
  assign memory[ 570 ] = 32'h00184463;
  assign memory[ 571 ] = 32'hFC32F7FF;
  assign memory[ 572 ] = 32'h2308E033;
  assign memory[ 573 ] = 32'h9B09930B;
  assign memory[ 574 ] = 32'h009222FA;
  assign memory[ 575 ] = 32'h9B0A435A;
  assign memory[ 576 ] = 32'h434B2164;
  assign memory[ 577 ] = 32'h9A0B18D1;
  assign memory[ 578 ] = 32'h009B0013;
  assign memory[ 579 ] = 32'h005B189B;
  assign memory[ 580 ] = 32'h9B0C18CA;
  assign memory[ 581 ] = 32'h228018D3;
  assign memory[ 582 ] = 32'h46940592;
  assign memory[ 583 ] = 32'h00184463;
  assign memory[ 584 ] = 32'hFC18F7FF;
  assign memory[ 585 ] = 32'h2309E019;
  assign memory[ 586 ] = 32'h9B09930B;
  assign memory[ 587 ] = 32'h009222FA;
  assign memory[ 588 ] = 32'h9B0A435A;
  assign memory[ 589 ] = 32'h434B2164;
  assign memory[ 590 ] = 32'h9A0B18D1;
  assign memory[ 591 ] = 32'h009B0013;
  assign memory[ 592 ] = 32'h005B189B;
  assign memory[ 593 ] = 32'h9B0C18CA;
  assign memory[ 594 ] = 32'h228018D3;
  assign memory[ 595 ] = 32'h46940592;
  assign memory[ 596 ] = 32'h00184463;
  assign memory[ 597 ] = 32'hFBFEF7FF;
  assign memory[ 598 ] = 32'hE2B446C0;
  assign memory[ 599 ] = 32'h2B099B10;
  assign memory[ 600 ] = 32'hE2B3D900;
  assign memory[ 601 ] = 32'h009A9B10;
  assign memory[ 602 ] = 32'h18D34B6A;
  assign memory[ 603 ] = 32'h469F681B;
  assign memory[ 604 ] = 32'h930A2300;
  assign memory[ 605 ] = 32'h22FA9B09;
  assign memory[ 606 ] = 32'h435A0092;
  assign memory[ 607 ] = 32'h21649B0A;
  assign memory[ 608 ] = 32'h18D1434B;
  assign memory[ 609 ] = 32'h00139A0B;
  assign memory[ 610 ] = 32'h189B009B;
  assign memory[ 611 ] = 32'h18CA005B;
  assign memory[ 612 ] = 32'h18D39B0C;
  assign memory[ 613 ] = 32'h05922280;
  assign memory[ 614 ] = 32'h44634694;
  assign memory[ 615 ] = 32'hF7FF0018;
  assign memory[ 616 ] = 32'hE0EDFBD9;
  assign memory[ 617 ] = 32'h930A2301;
  assign memory[ 618 ] = 32'h22FA9B09;
  assign memory[ 619 ] = 32'h435A0092;
  assign memory[ 620 ] = 32'h21649B0A;
  assign memory[ 621 ] = 32'h18D1434B;
  assign memory[ 622 ] = 32'h00139A0B;
  assign memory[ 623 ] = 32'h189B009B;
  assign memory[ 624 ] = 32'h18CA005B;
  assign memory[ 625 ] = 32'h18D39B0C;
  assign memory[ 626 ] = 32'h05922280;
  assign memory[ 627 ] = 32'h44634694;
  assign memory[ 628 ] = 32'hF7FF0018;
  assign memory[ 629 ] = 32'hE0D3FBBF;
  assign memory[ 630 ] = 32'h930A2302;
  assign memory[ 631 ] = 32'h22FA9B09;
  assign memory[ 632 ] = 32'h435A0092;
  assign memory[ 633 ] = 32'h21649B0A;
  assign memory[ 634 ] = 32'h18D1434B;
  assign memory[ 635 ] = 32'h00139A0B;
  assign memory[ 636 ] = 32'h189B009B;
  assign memory[ 637 ] = 32'h18CA005B;
  assign memory[ 638 ] = 32'h18D39B0C;
  assign memory[ 639 ] = 32'h05922280;
  assign memory[ 640 ] = 32'h44634694;
  assign memory[ 641 ] = 32'hF7FF0018;
  assign memory[ 642 ] = 32'hE0B9FBA5;
  assign memory[ 643 ] = 32'h930A2303;
  assign memory[ 644 ] = 32'h22FA9B09;
  assign memory[ 645 ] = 32'h435A0092;
  assign memory[ 646 ] = 32'h21649B0A;
  assign memory[ 647 ] = 32'h18D1434B;
  assign memory[ 648 ] = 32'h00139A0B;
  assign memory[ 649 ] = 32'h189B009B;
  assign memory[ 650 ] = 32'h18CA005B;
  assign memory[ 651 ] = 32'h18D39B0C;
  assign memory[ 652 ] = 32'h05922280;
  assign memory[ 653 ] = 32'h44634694;
  assign memory[ 654 ] = 32'hF7FF0018;
  assign memory[ 655 ] = 32'hE09FFB8B;
  assign memory[ 656 ] = 32'h930A2304;
  assign memory[ 657 ] = 32'h22FA9B09;
  assign memory[ 658 ] = 32'h435A0092;
  assign memory[ 659 ] = 32'h21649B0A;
  assign memory[ 660 ] = 32'h18D1434B;
  assign memory[ 661 ] = 32'h00139A0B;
  assign memory[ 662 ] = 32'h189B009B;
  assign memory[ 663 ] = 32'h18CA005B;
  assign memory[ 664 ] = 32'h18D39B0C;
  assign memory[ 665 ] = 32'h05922280;
  assign memory[ 666 ] = 32'h44634694;
  assign memory[ 667 ] = 32'hF7FF0018;
  assign memory[ 668 ] = 32'hE085FB71;
  assign memory[ 669 ] = 32'h930A2305;
  assign memory[ 670 ] = 32'h22FA9B09;
  assign memory[ 671 ] = 32'h435A0092;
  assign memory[ 672 ] = 32'h21649B0A;
  assign memory[ 673 ] = 32'h18D1434B;
  assign memory[ 674 ] = 32'h00139A0B;
  assign memory[ 675 ] = 32'h189B009B;
  assign memory[ 676 ] = 32'h18CA005B;
  assign memory[ 677 ] = 32'h18D39B0C;
  assign memory[ 678 ] = 32'h05922280;
  assign memory[ 679 ] = 32'h44634694;
  assign memory[ 680 ] = 32'hF7FF0018;
  assign memory[ 681 ] = 32'hE06BFB57;
  assign memory[ 682 ] = 32'h930A2306;
  assign memory[ 683 ] = 32'h22FA9B09;
  assign memory[ 684 ] = 32'h435A0092;
  assign memory[ 685 ] = 32'h21649B0A;
  assign memory[ 686 ] = 32'h18D1434B;
  assign memory[ 687 ] = 32'h00139A0B;
  assign memory[ 688 ] = 32'h189B009B;
  assign memory[ 689 ] = 32'h18CA005B;
  assign memory[ 690 ] = 32'h18D39B0C;
  assign memory[ 691 ] = 32'h05922280;
  assign memory[ 692 ] = 32'h44634694;
  assign memory[ 693 ] = 32'hF7FF0018;
  assign memory[ 694 ] = 32'hE051FB3D;
  assign memory[ 695 ] = 32'h930A2307;
  assign memory[ 696 ] = 32'h22FA9B09;
  assign memory[ 697 ] = 32'h435A0092;
  assign memory[ 698 ] = 32'h21649B0A;
  assign memory[ 699 ] = 32'h18D1434B;
  assign memory[ 700 ] = 32'h00139A0B;
  assign memory[ 701 ] = 32'h189B009B;
  assign memory[ 702 ] = 32'h18CA005B;
  assign memory[ 703 ] = 32'h18D39B0C;
  assign memory[ 704 ] = 32'h05922280;
  assign memory[ 705 ] = 32'h44634694;
  assign memory[ 706 ] = 32'hF7FF0018;
  assign memory[ 707 ] = 32'hE037FB23;
  assign memory[ 708 ] = 32'h000010E8;
  assign memory[ 709 ] = 32'h00001110;
  assign memory[ 710 ] = 32'h930A2308;
  assign memory[ 711 ] = 32'h22FA9B09;
  assign memory[ 712 ] = 32'h435A0092;
  assign memory[ 713 ] = 32'h21649B0A;
  assign memory[ 714 ] = 32'h18D1434B;
  assign memory[ 715 ] = 32'h00139A0B;
  assign memory[ 716 ] = 32'h189B009B;
  assign memory[ 717 ] = 32'h18CA005B;
  assign memory[ 718 ] = 32'h18D39B0C;
  assign memory[ 719 ] = 32'h05922280;
  assign memory[ 720 ] = 32'h44634694;
  assign memory[ 721 ] = 32'hF7FF0018;
  assign memory[ 722 ] = 32'hE019FB05;
  assign memory[ 723 ] = 32'h930A2309;
  assign memory[ 724 ] = 32'h22FA9B09;
  assign memory[ 725 ] = 32'h435A0092;
  assign memory[ 726 ] = 32'h21649B0A;
  assign memory[ 727 ] = 32'h18D1434B;
  assign memory[ 728 ] = 32'h00139A0B;
  assign memory[ 729 ] = 32'h189B009B;
  assign memory[ 730 ] = 32'h18CA005B;
  assign memory[ 731 ] = 32'h18D39B0C;
  assign memory[ 732 ] = 32'h05922280;
  assign memory[ 733 ] = 32'h44634694;
  assign memory[ 734 ] = 32'hF7FF0018;
  assign memory[ 735 ] = 32'h46C0FAEB;
  assign memory[ 736 ] = 32'h9B10E1A4;
  assign memory[ 737 ] = 32'hD9002B09;
  assign memory[ 738 ] = 32'h9B10E1A3;
  assign memory[ 739 ] = 32'h4BD2009A;
  assign memory[ 740 ] = 32'h681B18D3;
  assign memory[ 741 ] = 32'h2300469F;
  assign memory[ 742 ] = 32'h9B099309;
  assign memory[ 743 ] = 32'h009222FA;
  assign memory[ 744 ] = 32'h9B0A435A;
  assign memory[ 745 ] = 32'h434B2164;
  assign memory[ 746 ] = 32'h9A0B18D1;
  assign memory[ 747 ] = 32'h009B0013;
  assign memory[ 748 ] = 32'h005B189B;
  assign memory[ 749 ] = 32'h9B0C18CA;
  assign memory[ 750 ] = 32'h228018D3;
  assign memory[ 751 ] = 32'h46940592;
  assign memory[ 752 ] = 32'h00184463;
  assign memory[ 753 ] = 32'hFAC6F7FF;
  assign memory[ 754 ] = 32'h2301E0E9;
  assign memory[ 755 ] = 32'h9B099309;
  assign memory[ 756 ] = 32'h009222FA;
  assign memory[ 757 ] = 32'h9B0A435A;
  assign memory[ 758 ] = 32'h434B2164;
  assign memory[ 759 ] = 32'h9A0B18D1;
  assign memory[ 760 ] = 32'h009B0013;
  assign memory[ 761 ] = 32'h005B189B;
  assign memory[ 762 ] = 32'h9B0C18CA;
  assign memory[ 763 ] = 32'h228018D3;
  assign memory[ 764 ] = 32'h46940592;
  assign memory[ 765 ] = 32'h00184463;
  assign memory[ 766 ] = 32'hFAACF7FF;
  assign memory[ 767 ] = 32'h2302E0CF;
  assign memory[ 768 ] = 32'h9B099309;
  assign memory[ 769 ] = 32'h009222FA;
  assign memory[ 770 ] = 32'h9B0A435A;
  assign memory[ 771 ] = 32'h434B2164;
  assign memory[ 772 ] = 32'h9A0B18D1;
  assign memory[ 773 ] = 32'h009B0013;
  assign memory[ 774 ] = 32'h005B189B;
  assign memory[ 775 ] = 32'h9B0C18CA;
  assign memory[ 776 ] = 32'h228018D3;
  assign memory[ 777 ] = 32'h46940592;
  assign memory[ 778 ] = 32'h00184463;
  assign memory[ 779 ] = 32'hFA92F7FF;
  assign memory[ 780 ] = 32'h2303E0B5;
  assign memory[ 781 ] = 32'h9B099309;
  assign memory[ 782 ] = 32'h009222FA;
  assign memory[ 783 ] = 32'h9B0A435A;
  assign memory[ 784 ] = 32'h434B2164;
  assign memory[ 785 ] = 32'h9A0B18D1;
  assign memory[ 786 ] = 32'h009B0013;
  assign memory[ 787 ] = 32'h005B189B;
  assign memory[ 788 ] = 32'h9B0C18CA;
  assign memory[ 789 ] = 32'h228018D3;
  assign memory[ 790 ] = 32'h46940592;
  assign memory[ 791 ] = 32'h00184463;
  assign memory[ 792 ] = 32'hFA78F7FF;
  assign memory[ 793 ] = 32'h2304E09B;
  assign memory[ 794 ] = 32'h9B099309;
  assign memory[ 795 ] = 32'h009222FA;
  assign memory[ 796 ] = 32'h9B0A435A;
  assign memory[ 797 ] = 32'h434B2164;
  assign memory[ 798 ] = 32'h9A0B18D1;
  assign memory[ 799 ] = 32'h009B0013;
  assign memory[ 800 ] = 32'h005B189B;
  assign memory[ 801 ] = 32'h9B0C18CA;
  assign memory[ 802 ] = 32'h228018D3;
  assign memory[ 803 ] = 32'h46940592;
  assign memory[ 804 ] = 32'h00184463;
  assign memory[ 805 ] = 32'hFA5EF7FF;
  assign memory[ 806 ] = 32'h2305E081;
  assign memory[ 807 ] = 32'h9B099309;
  assign memory[ 808 ] = 32'h009222FA;
  assign memory[ 809 ] = 32'h9B0A435A;
  assign memory[ 810 ] = 32'h434B2164;
  assign memory[ 811 ] = 32'h9A0B18D1;
  assign memory[ 812 ] = 32'h009B0013;
  assign memory[ 813 ] = 32'h005B189B;
  assign memory[ 814 ] = 32'h9B0C18CA;
  assign memory[ 815 ] = 32'h228018D3;
  assign memory[ 816 ] = 32'h46940592;
  assign memory[ 817 ] = 32'h00184463;
  assign memory[ 818 ] = 32'hFA44F7FF;
  assign memory[ 819 ] = 32'h2306E067;
  assign memory[ 820 ] = 32'h9B099309;
  assign memory[ 821 ] = 32'h009222FA;
  assign memory[ 822 ] = 32'h9B0A435A;
  assign memory[ 823 ] = 32'h434B2164;
  assign memory[ 824 ] = 32'h9A0B18D1;
  assign memory[ 825 ] = 32'h009B0013;
  assign memory[ 826 ] = 32'h005B189B;
  assign memory[ 827 ] = 32'h9B0C18CA;
  assign memory[ 828 ] = 32'h228018D3;
  assign memory[ 829 ] = 32'h46940592;
  assign memory[ 830 ] = 32'h00184463;
  assign memory[ 831 ] = 32'hFA2AF7FF;
  assign memory[ 832 ] = 32'h2307E04D;
  assign memory[ 833 ] = 32'h9B099309;
  assign memory[ 834 ] = 32'h009222FA;
  assign memory[ 835 ] = 32'h9B0A435A;
  assign memory[ 836 ] = 32'h434B2164;
  assign memory[ 837 ] = 32'h9A0B18D1;
  assign memory[ 838 ] = 32'h009B0013;
  assign memory[ 839 ] = 32'h005B189B;
  assign memory[ 840 ] = 32'h9B0C18CA;
  assign memory[ 841 ] = 32'h228018D3;
  assign memory[ 842 ] = 32'h46940592;
  assign memory[ 843 ] = 32'h00184463;
  assign memory[ 844 ] = 32'hFA10F7FF;
  assign memory[ 845 ] = 32'h2308E033;
  assign memory[ 846 ] = 32'h9B099309;
  assign memory[ 847 ] = 32'h009222FA;
  assign memory[ 848 ] = 32'h9B0A435A;
  assign memory[ 849 ] = 32'h434B2164;
  assign memory[ 850 ] = 32'h9A0B18D1;
  assign memory[ 851 ] = 32'h009B0013;
  assign memory[ 852 ] = 32'h005B189B;
  assign memory[ 853 ] = 32'h9B0C18CA;
  assign memory[ 854 ] = 32'h228018D3;
  assign memory[ 855 ] = 32'h46940592;
  assign memory[ 856 ] = 32'h00184463;
  assign memory[ 857 ] = 32'hF9F6F7FF;
  assign memory[ 858 ] = 32'h2309E019;
  assign memory[ 859 ] = 32'h9B099309;
  assign memory[ 860 ] = 32'h009222FA;
  assign memory[ 861 ] = 32'h9B0A435A;
  assign memory[ 862 ] = 32'h434B2164;
  assign memory[ 863 ] = 32'h9A0B18D1;
  assign memory[ 864 ] = 32'h009B0013;
  assign memory[ 865 ] = 32'h005B189B;
  assign memory[ 866 ] = 32'h9B0C18CA;
  assign memory[ 867 ] = 32'h228018D3;
  assign memory[ 868 ] = 32'h46940592;
  assign memory[ 869 ] = 32'h00184463;
  assign memory[ 870 ] = 32'hF9DCF7FF;
  assign memory[ 871 ] = 32'h46C046C0;
  assign memory[ 872 ] = 32'h9A07E097;
  assign memory[ 873 ] = 32'h33FF2340;
  assign memory[ 874 ] = 32'hDD04429A;
  assign memory[ 875 ] = 32'h2B009B08;
  assign memory[ 876 ] = 32'h2301D101;
  assign memory[ 877 ] = 32'h9B07930F;
  assign memory[ 878 ] = 32'hD1122B00;
  assign memory[ 879 ] = 32'h2B019B0F;
  assign memory[ 880 ] = 32'h9B08D10F;
  assign memory[ 881 ] = 32'hD10C2B00;
  assign memory[ 882 ] = 32'h2B049B15;
  assign memory[ 883 ] = 32'h9B15DC05;
  assign memory[ 884 ] = 32'h93153301;
  assign memory[ 885 ] = 32'h930F2300;
  assign memory[ 886 ] = 32'h2300E003;
  assign memory[ 887 ] = 32'h23009315;
  assign memory[ 888 ] = 32'h9B15930F;
  assign memory[ 889 ] = 32'hD9012B05;
  assign memory[ 890 ] = 32'hFAC8F7FF;
  assign memory[ 891 ] = 32'h009A9B15;
  assign memory[ 892 ] = 32'h18D34B3A;
  assign memory[ 893 ] = 32'h469F681B;
  assign memory[ 894 ] = 32'hF7FF2002;
  assign memory[ 895 ] = 32'h0003F9C3;
  assign memory[ 896 ] = 32'h9A139306;
  assign memory[ 897 ] = 32'h00119B06;
  assign memory[ 898 ] = 32'hF7FF0018;
  assign memory[ 899 ] = 32'h0003F9DF;
  assign memory[ 900 ] = 32'hF7FF0018;
  assign memory[ 901 ] = 32'hE05DF99F;
  assign memory[ 902 ] = 32'hF7FF2003;
  assign memory[ 903 ] = 32'h0003F9B3;
  assign memory[ 904 ] = 32'h9B059305;
  assign memory[ 905 ] = 32'hF7FF0018;
  assign memory[ 906 ] = 32'h0003F9EF;
  assign memory[ 907 ] = 32'hF7FF0018;
  assign memory[ 908 ] = 32'hE04FF991;
  assign memory[ 909 ] = 32'hF7FF2004;
  assign memory[ 910 ] = 32'h0003F9A5;
  assign memory[ 911 ] = 32'h9B049304;
  assign memory[ 912 ] = 32'hF7FF0018;
  assign memory[ 913 ] = 32'h0003FA0D;
  assign memory[ 914 ] = 32'hF7FF0018;
  assign memory[ 915 ] = 32'hE041F983;
  assign memory[ 916 ] = 32'h00189B02;
  assign memory[ 917 ] = 32'hF97EF7FF;
  assign memory[ 918 ] = 32'h9B12E03C;
  assign memory[ 919 ] = 32'h061222C0;
  assign memory[ 920 ] = 32'h44634694;
  assign memory[ 921 ] = 32'hF7FF0018;
  assign memory[ 922 ] = 32'hE033F975;
  assign memory[ 923 ] = 32'hF7FF2002;
  assign memory[ 924 ] = 32'h0003F989;
  assign memory[ 925 ] = 32'h20039306;
  assign memory[ 926 ] = 32'hF984F7FF;
  assign memory[ 927 ] = 32'h93050003;
  assign memory[ 928 ] = 32'h9A139B06;
  assign memory[ 929 ] = 32'h0013435A;
  assign memory[ 930 ] = 32'h189B009B;
  assign memory[ 931 ] = 32'h4914005B;
  assign memory[ 932 ] = 32'hF0000018;
  assign memory[ 933 ] = 32'h0003F829;
  assign memory[ 934 ] = 32'h9B05001C;
  assign memory[ 935 ] = 32'h00184911;
  assign memory[ 936 ] = 32'hF822F000;
  assign memory[ 937 ] = 32'h00190003;
  assign memory[ 938 ] = 32'hF0000020;
  assign memory[ 939 ] = 32'h0003F81D;
  assign memory[ 940 ] = 32'h061222E0;
  assign memory[ 941 ] = 32'h44634694;
  assign memory[ 942 ] = 32'hF7FF0018;
  assign memory[ 943 ] = 32'hE009F94B;
  assign memory[ 944 ] = 32'hF7FF46C0;
  assign memory[ 945 ] = 32'h46C0FA5B;
  assign memory[ 946 ] = 32'hFA58F7FF;
  assign memory[ 947 ] = 32'hF7FF46C0;
  assign memory[ 948 ] = 32'h46C0FA55;
  assign memory[ 949 ] = 32'hFA52F7FF;
  assign memory[ 950 ] = 32'h00001138;
  assign memory[ 951 ] = 32'h00001160;
  assign memory[ 952 ] = 32'h000F4240;
  assign memory[ 953 ] = 32'h02BF2000;
  assign memory[ 954 ] = 32'h430B4603;
  assign memory[ 955 ] = 32'h2200D47F;
  assign memory[ 956 ] = 32'h428B0843;
  assign memory[ 957 ] = 32'h0903D374;
  assign memory[ 958 ] = 32'hD35F428B;
  assign memory[ 959 ] = 32'h428B0A03;
  assign memory[ 960 ] = 32'h0B03D344;
  assign memory[ 961 ] = 32'hD328428B;
  assign memory[ 962 ] = 32'h428B0C03;
  assign memory[ 963 ] = 32'h22FFD30D;
  assign memory[ 964 ] = 32'hBA120209;
  assign memory[ 965 ] = 32'h428B0C03;
  assign memory[ 966 ] = 32'h1212D302;
  assign memory[ 967 ] = 32'hD0650209;
  assign memory[ 968 ] = 32'h428B0B03;
  assign memory[ 969 ] = 32'hE000D319;
  assign memory[ 970 ] = 32'h0BC30A09;
  assign memory[ 971 ] = 32'hD301428B;
  assign memory[ 972 ] = 32'h1AC003CB;
  assign memory[ 973 ] = 32'h0B834152;
  assign memory[ 974 ] = 32'hD301428B;
  assign memory[ 975 ] = 32'h1AC0038B;
  assign memory[ 976 ] = 32'h0B434152;
  assign memory[ 977 ] = 32'hD301428B;
  assign memory[ 978 ] = 32'h1AC0034B;
  assign memory[ 979 ] = 32'h0B034152;
  assign memory[ 980 ] = 32'hD301428B;
  assign memory[ 981 ] = 32'h1AC0030B;
  assign memory[ 982 ] = 32'h0AC34152;
  assign memory[ 983 ] = 32'hD301428B;
  assign memory[ 984 ] = 32'h1AC002CB;
  assign memory[ 985 ] = 32'h0A834152;
  assign memory[ 986 ] = 32'hD301428B;
  assign memory[ 987 ] = 32'h1AC0028B;
  assign memory[ 988 ] = 32'h0A434152;
  assign memory[ 989 ] = 32'hD301428B;
  assign memory[ 990 ] = 32'h1AC0024B;
  assign memory[ 991 ] = 32'h0A034152;
  assign memory[ 992 ] = 32'hD301428B;
  assign memory[ 993 ] = 32'h1AC0020B;
  assign memory[ 994 ] = 32'hD2CD4152;
  assign memory[ 995 ] = 32'h428B09C3;
  assign memory[ 996 ] = 32'h01CBD301;
  assign memory[ 997 ] = 32'h41521AC0;
  assign memory[ 998 ] = 32'h428B0983;
  assign memory[ 999 ] = 32'h018BD301;
  assign memory[ 1000 ] = 32'h41521AC0;
  assign memory[ 1001 ] = 32'h428B0943;
  assign memory[ 1002 ] = 32'h014BD301;
  assign memory[ 1003 ] = 32'h41521AC0;
  assign memory[ 1004 ] = 32'h428B0903;
  assign memory[ 1005 ] = 32'h010BD301;
  assign memory[ 1006 ] = 32'h41521AC0;
  assign memory[ 1007 ] = 32'h428B08C3;
  assign memory[ 1008 ] = 32'h00CBD301;
  assign memory[ 1009 ] = 32'h41521AC0;
  assign memory[ 1010 ] = 32'h428B0883;
  assign memory[ 1011 ] = 32'h008BD301;
  assign memory[ 1012 ] = 32'h41521AC0;
  assign memory[ 1013 ] = 32'h428B0843;
  assign memory[ 1014 ] = 32'h004BD301;
  assign memory[ 1015 ] = 32'h41521AC0;
  assign memory[ 1016 ] = 32'hD2001A41;
  assign memory[ 1017 ] = 32'h41524601;
  assign memory[ 1018 ] = 32'h47704610;
  assign memory[ 1019 ] = 32'h0FCAE05D;
  assign memory[ 1020 ] = 32'h4249D000;
  assign memory[ 1021 ] = 32'hD3001003;
  assign memory[ 1022 ] = 32'h40534240;
  assign memory[ 1023 ] = 32'h469C2200;
  assign memory[ 1024 ] = 32'h428B0903;
  assign memory[ 1025 ] = 32'h0A03D32D;
  assign memory[ 1026 ] = 32'hD312428B;
  assign memory[ 1027 ] = 32'h018922FC;
  assign memory[ 1028 ] = 32'h0A03BA12;
  assign memory[ 1029 ] = 32'hD30C428B;
  assign memory[ 1030 ] = 32'h11920189;
  assign memory[ 1031 ] = 32'hD308428B;
  assign memory[ 1032 ] = 32'h11920189;
  assign memory[ 1033 ] = 32'hD304428B;
  assign memory[ 1034 ] = 32'hD03A0189;
  assign memory[ 1035 ] = 32'hE0001192;
  assign memory[ 1036 ] = 32'h09C30989;
  assign memory[ 1037 ] = 32'hD301428B;
  assign memory[ 1038 ] = 32'h1AC001CB;
  assign memory[ 1039 ] = 32'h09834152;
  assign memory[ 1040 ] = 32'hD301428B;
  assign memory[ 1041 ] = 32'h1AC0018B;
  assign memory[ 1042 ] = 32'h09434152;
  assign memory[ 1043 ] = 32'hD301428B;
  assign memory[ 1044 ] = 32'h1AC0014B;
  assign memory[ 1045 ] = 32'h09034152;
  assign memory[ 1046 ] = 32'hD301428B;
  assign memory[ 1047 ] = 32'h1AC0010B;
  assign memory[ 1048 ] = 32'h08C34152;
  assign memory[ 1049 ] = 32'hD301428B;
  assign memory[ 1050 ] = 32'h1AC000CB;
  assign memory[ 1051 ] = 32'h08834152;
  assign memory[ 1052 ] = 32'hD301428B;
  assign memory[ 1053 ] = 32'h1AC0008B;
  assign memory[ 1054 ] = 32'hD2D94152;
  assign memory[ 1055 ] = 32'h428B0843;
  assign memory[ 1056 ] = 32'h004BD301;
  assign memory[ 1057 ] = 32'h41521AC0;
  assign memory[ 1058 ] = 32'hD2001A41;
  assign memory[ 1059 ] = 32'h46634601;
  assign memory[ 1060 ] = 32'h105B4152;
  assign memory[ 1061 ] = 32'hD3014610;
  assign memory[ 1062 ] = 32'h2B004240;
  assign memory[ 1063 ] = 32'h4249D500;
  assign memory[ 1064 ] = 32'h46634770;
  assign memory[ 1065 ] = 32'hD300105B;
  assign memory[ 1066 ] = 32'hB5014240;
  assign memory[ 1067 ] = 32'hF0002000;
  assign memory[ 1068 ] = 32'hBD02F805;
  assign memory[ 1069 ] = 32'hD0F82900;
  assign memory[ 1070 ] = 32'h4770E716;
  assign memory[ 1071 ] = 32'h46C04770;
  assign memory[ 1072 ] = 32'h00000528;
  assign memory[ 1073 ] = 32'h0000055C;
  assign memory[ 1074 ] = 32'h00000590;
  assign memory[ 1075 ] = 32'h000005C4;
  assign memory[ 1076 ] = 32'h000005F8;
  assign memory[ 1077 ] = 32'h0000062C;
  assign memory[ 1078 ] = 32'h00000660;
  assign memory[ 1079 ] = 32'h00000694;
  assign memory[ 1080 ] = 32'h000006D4;
  assign memory[ 1081 ] = 32'h00000708;
  assign memory[ 1082 ] = 32'h00000752;
  assign memory[ 1083 ] = 32'h00000786;
  assign memory[ 1084 ] = 32'h000007BA;
  assign memory[ 1085 ] = 32'h000007EE;
  assign memory[ 1086 ] = 32'h00000822;
  assign memory[ 1087 ] = 32'h00000856;
  assign memory[ 1088 ] = 32'h0000088A;
  assign memory[ 1089 ] = 32'h000008BE;
  assign memory[ 1090 ] = 32'h000008F2;
  assign memory[ 1091 ] = 32'h00000926;
  assign memory[ 1092 ] = 32'h00000970;
  assign memory[ 1093 ] = 32'h000009A4;
  assign memory[ 1094 ] = 32'h000009D8;
  assign memory[ 1095 ] = 32'h00000A0C;
  assign memory[ 1096 ] = 32'h00000A40;
  assign memory[ 1097 ] = 32'h00000A74;
  assign memory[ 1098 ] = 32'h00000AA8;
  assign memory[ 1099 ] = 32'h00000ADC;
  assign memory[ 1100 ] = 32'h00000B18;
  assign memory[ 1101 ] = 32'h00000B4C;
  assign memory[ 1102 ] = 32'h00000B96;
  assign memory[ 1103 ] = 32'h00000BCA;
  assign memory[ 1104 ] = 32'h00000BFE;
  assign memory[ 1105 ] = 32'h00000C32;
  assign memory[ 1106 ] = 32'h00000C66;
  assign memory[ 1107 ] = 32'h00000C9A;
  assign memory[ 1108 ] = 32'h00000CCE;
  assign memory[ 1109 ] = 32'h00000D02;
  assign memory[ 1110 ] = 32'h00000D36;
  assign memory[ 1111 ] = 32'h00000D6A;
  assign memory[ 1112 ] = 32'h00000DF8;
  assign memory[ 1113 ] = 32'h00000E18;
  assign memory[ 1114 ] = 32'h00000E34;
  assign memory[ 1115 ] = 32'h00000E50;
  assign memory[ 1116 ] = 32'h00000E5A;
  assign memory[ 1117 ] = 32'h00000E6C;
  assign memory[ 1118 ] = 32'h40000000;
  assign memory[ 1119 ] = 32'h50000000;
//Generate the control signals in the address phase
  always_ff @(posedge HCLK, negedge HRESETn)
    if (! HRESETn )
      begin
        read_enable <= '0;
        word_address <= '0;
        byte_select <= '0;
      end
    else if ( HREADY && HSEL && (HTRANS != No_Transfer) )
      begin
        read_enable <= ! HWRITE;
        word_address <= HADDR[MEMWIDTH:2];
        byte_select <= generate_byte_select( HSIZE, HADDR[1:0] );
     end
    else
      begin
        read_enable <= '0;
        word_address <= '0;
        byte_select <= '0;
     end

//Act on control signals in the data phase

  // no write since thisis a ROM

  //read
  // (output of zero when not enabled for read is not necessary but may help with debugging)
  assign HRDATA[ 7: 0] = ( read_enable && byte_select[0] ) ? memory[word_address][ 7: 0] : '0;
  assign HRDATA[15: 8] = ( read_enable && byte_select[1] ) ? memory[word_address][15: 8] : '0;
  assign HRDATA[23:16] = ( read_enable && byte_select[2] ) ? memory[word_address][23:16] : '0;
  assign HRDATA[31:24] = ( read_enable && byte_select[3] ) ? memory[word_address][31:24] : '0;

//Transfer Response
  assign HREADYOUT = '1; //Single cycle Write & Read. Zero Wait state operations


// decode byte select signals from the size and the lowest two address bits
  function logic [3:0] generate_byte_select( logic [2:0] size, logic [1:0] byte_adress );
    logic byte3, byte2, byte1, byte0;
    byte0 = size[1] || ( byte_adress == 0 );
    byte1 = size[1] || ( size[0] && ( byte_adress == 0 ) ) || ( byte_adress == 1 );
    byte2 = size[1] || ( byte_adress == 2 );
    byte3 = size[1] || ( size[0] && ( byte_adress == 2 ) ) || ( byte_adress == 3 );
    return { byte3, byte2, byte1, byte0 };
  endfunction

endmodule

